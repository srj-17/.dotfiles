library IEEE;
use IEEE.std_logic_1164.all

entity andGate is
    port(A: in std_logic